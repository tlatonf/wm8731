// Copyright (c) 2024 Tlatonf

`define NO_TAPS         100
`define WIDTH_DATA      24
`define WIDTH_COEFF     20


`define WIDTH_PROC      `WIDTH_DATA + `WIDTH_COEFF
`define WIDTH_SUM       `WIDTH_PROC + 1

`define FILE_COEFF      "coefficient.bin"

//`define FILE_TB_INPUT   "../10_material/sine.hex"
//`define FILE_TB_OUTPUT  "../10_material/output.hex"
